module full_adder_1bit_LS_series(A, B, Carry_in, SUM, Carry_out);
  input A;
  input B;
  input Carry_in;
  output SUM;
  output Carry_out;

  wire x;
  wire y;
  wire z;

  IC74LS86 xor_ic_inst( ...complete the code in lab ...
  IC74LS08 and_ic_inst( ...complete the code in lab ...
  IC74LS32 or_ic_inst( ...complete the code in lab ...

endmodule